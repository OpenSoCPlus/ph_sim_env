/*====================================

     MODULE : @TOP_MODULE@
     AUTHOR : @AUTHOR@

====================================*/
module @TOP_MODULE@(
	rstn      ,
	clk        
);


//=====================================
//
//          PARAMETERS 
//
//=====================================


//=====================================
//
//          I/O PORTS 
//
//=====================================
input        rstn      ; 
input        clk       ;

//=====================================
//
//          REGISTERS
//
//=====================================


//=====================================
//
//          WIRES
//
//=====================================


//=====================================
//
//          MAIN
//
//=====================================


endmodule


